module Test(
input a, 
input b, 
input c,
output l1,
output l2, 
output l3
);

assign l1 = a;
assign l2 = b;
assign l3 = c;

endmodule